`timescale 1ns/1ps

module user_def;
	defparam soc_tb.m_uart.Input_Udata = "./inputs/soc_top/sim/tests/s_1_261_bb_rom_cmd_sleep_hw_adv_has_sleep/uart.cm";
endmodule
