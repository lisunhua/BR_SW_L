`timescale 1ns/1ps

module user_def;
	//defparam  u_agc_sim_m.IQ_DATA_PATH = "./inputs/soc_top/sim/tests/s_1_2A3_bb_bt_le_agc_dtm_1m_rx/iq_data_ble_1m_tx.txt";
endmodule
