`timescale 1ns/1ps


module user_def;
	defparam  u_pcm_sim.PCM_DATA_PATH = "./inputs/soc_top/sim/tests/d_1_240_bb_bt_br_2-ev3_pcm55/sine_snd_data.txt";
endmodule
