`timescale 1ns/1ps

module user_def;
	defparam  CLT.u_spi_flash0.Init_File = "./inputs/soc_top/sim/tests/d_1_002_scu_remap_flash/flash_clt.hex";
	defparam  SVR.u_spi_flash0.Init_File = "./inputs/soc_top/sim/tests/d_1_002_scu_remap_flash/flash_svr.hex";
endmodule
