//Automatically generate file.

`include "inputs/soc_top/sim/tb/inc/chip_def.inc"

   reg [6:0] error_count;

task ana_connect_dig;

//===========================================
   error_count = 0;

   for (int i=0; i<40; i++) begin

    #100;
	force  `IOMUX_XRM.scan_test_clock  = $urandom;
	force  `PAD_XRM.u_TEST_PAD.C = $urandom;
	force  `IOMUX_XRM.scan_test_clock = $urandom;
	force  `PAD_XRM.u_TEST_PAD.C = $urandom;
	force  `IOMUX_XRM.sw_test_en = $urandom;
	force  `IOMUX_XRM.rf_test_en = $urandom;
	force  `IOMUX_XRM.bb_test_en = $urandom;
	force  `IOMUX_XRM.mbist_test_en = $urandom;
	force  `IOMUX_XRM.bsd_test_en = $urandom;
	force  `ANA_XRM.CLK_26M_OUT = $urandom;
	force  `CLK_XRM.clk_24m_rf = $urandom;
	force  `ANA_XRM.ADC_DATA[10:0] = $urandom;
	force  `ANA_XRM.ADC_VDET_INDEX = $urandom;
	force  `ANA_XRM.DCDC_OCP_DET = $urandom;
	force  `ANA_XRM.DCDC_PWM_TEST = $urandom;
	force  `ANA_XRM.DCDC_START_TEST = $urandom;
	force  `ANA_XRM.DCDC_ZCD_TEST = $urandom;
	force  `ANA_XRM.DPLL_LOCK = $urandom;
	force  `ANA_XRM.DPLL_OUT_16M = $urandom;
	force  `ANA_XRM.DPLL_OUT_24M = $urandom;
	force  `ANA_XRM.DPLL_OUT_192M = $urandom;
	force  `ANA_XRM.DPLL_OUT_192M_TEST = $urandom;
	force  `ANA_XRM.LVD_BB = $urandom;
	force  `ANA_XRM.POR_BB = $urandom;
	force  `ANA_XRM.RCO32_CAL_CODE[13:0] = $urandom;
	force  `ANA_XRM.RCO32_COARSE_DONE = $urandom;
	force  `ANA_XRM.RCO32_FINE_DONE = $urandom;
	force  `ANA_XRM.RCO_32K_BB = $urandom;
	force  `SCU_XRM.ana_ctl4[11:10] = $urandom;
	force  `PAD_XRM.ADC_IN[3:0] = $urandom;
	force  `SCU_XRM.ana_ctl3[5:4] = $urandom;
	force  `SCU_XRM.ana_ctl3[8:6] = $urandom;
	force  `SCU_XRM.ana_ctl3[3] = $urandom;
	force  `SCU_XRM.ana_ctl3[2:0] = $urandom;
	force  `SCU_XRM.ana_ctl4[2] = $urandom;
	force  `SCU_XRM.ana_ctl4[1] = $urandom;
	force  `SCU_XRM.ana_ctl4[0] = $urandom;
	force  `SCU_XRM.ana_ctl4[12] = $urandom;
	force  `SCU_XRM.ana_ctl4[8:7] = $urandom;
	force  `SCU_XRM.ana_ctl4[6] = $urandom;
	force  `SCU_XRM.ana_ctl4[14:13] = $urandom;
	force  `SCU_XRM.ana_ctl4[18:15] = $urandom;
	force  `SCU_XRM.ana_ctl4[20:19] = $urandom;
	force  `SCU_XRM.ana_ctl0[12] = $urandom;
	force  `SCU_XRM.ana_ctl0[31] = $urandom;
	force  `SCU_XRM.ana_ctl0[29] = $urandom;
	force  `SCU_XRM.ana_ctl0[30] = $urandom;
	force  `SCU_XRM.ana_ctl0[22] = $urandom;
	force  `SCU_XRM.ana_ctl4[9] = $urandom;
	force  `CORE_XRM.bb_dac_i[10:0] = $urandom;
	force  `CORE_XRM.bb_dac_q[10:0] = $urandom;
	force   `CORE_XRM.bb_tx_gain[2:0] = $urandom;
	force  `SCUREG_XRM.ana_ctl2[29:16] = $urandom;
	force  `SCU_XRM.ana_ctl2[4:3] = $urandom;
	force  `SCUREG_XRM.ana_ctl2[14:13] = $urandom;
	force  `SCU_XRM.ana_ctl3[28:27] = $urandom;
	force  `SCU_XRM.ana_ctl1[18:16] = $urandom;
	force  `SCU_XRM.ana_ctl4[28:26] = $urandom;
	force  `SCU_XRM.ana_ctl4[23:21] = $urandom;
	force  `SCU_XRM.ana_ctl3[31:29] = $urandom;
	force  `SCU_XRM.ana_ctl1[4:2] = $urandom;
	force  `SCU_XRM.ana_ctl4[31:29] = $urandom;
	force  `SCU_XRM.ana_ctl4[5:3] = $urandom;
	force  `SCU_XRM.ana_ctl3[26:23] = $urandom;
	force  `SCU_XRM.ana_ctl1[12:7] = $urandom;
	force  `CORE_XRM.bb_freq_hop[6:0] = $urandom;
	force  `CORE_XRM.bb_rx_agc[7:0] = $urandom;
	force  `CORE_XRM.bb_temp_comp_tx_gain[7:0] = $urandom;
	force  `CLK_XRM.rf_adc_clk = $urandom;
	force  `CLK_XRM.clk_48m_bb = $urandom;
	force  `CORE_XRM.DA_RX_PKD_RSTN = $urandom;
	force  `SCU_XRM.ana_ctl0[4] = $urandom;
	force  `IOMUX_XRM.clk_ext_in = $urandom;
	force  `SCUREG_XRM.ana_ctl0[11] = $urandom;
	force  `SCUREG_XRM.ana_ctl0[19] = $urandom;
	force  `DUT_XRM.u_pad_ring.EN_CHIP_V33 = $urandom;
	force  `SCUREG_XRM.ana_ctl0[28] = $urandom;
	force  `SCUREG_XRM.ana_ctl0[15] = $urandom;
	force  `SCUREG_XRM.ana_ctl0[14] = $urandom;
	force  `SCUREG_XRM.ana_ctl0[17] = $urandom;
	force  `CLK_XRM.mux_dpll_sel = $urandom;
	force  `SCUREG_XRM.ana_ctl0[13] = $urandom;
	force  `SCUREG_XRM.ana_ctl0[25] = $urandom;
	force  `SCUREG_XRM.ana_ctl0[27] = $urandom;
	force  `CLK_XRM.mux_ldoxo_sel = $urandom;
	force  `SCUREG_XRM.ana_ctl1[23] = $urandom;
	force  `SCUREG_XRM.ana_ctl0[21] = $urandom;
	force  `SCUREG_XRM.ana_ctl0[18] = $urandom;
	force  `SCUREG_XRM.ana_ctl0[16] = $urandom;
	force  `SCUREG_XRM.ana_ctl1[5] = $urandom;
	force  `SCUREG_XRM.ana_ctl1[6] = $urandom;
	force  `SCUREG_XRM.ana_ctl1[15] = $urandom;
	force  `SCUREG_XRM.ana_ctl1[0] = $urandom;
	force  `SCUREG_XRM.ana_ctl1[1] = $urandom;
	force  `SCUREG_XRM.ana_ctl1[22] = $urandom;
	force  `SCUREG_XRM.ana_ctl2[31] = $urandom;
	force  `SCUREG_XRM.ana_ctl2[30] = $urandom;
	force  `SCUREG_XRM.ana_ctl2[15] = $urandom;
	force  `SCUREG_XRM.ana_ctl2[12] = $urandom;
	force  `IOMUX_XRM.resetn_rf = $urandom;
	force  `IOMUX_XRM.rf_spis_clk_ana = $urandom;
	force  `IOMUX_XRM.rf_spis_csn_ana = $urandom;
	force  `IOMUX_XRM.rf_spis_mosi_ana = $urandom;
	force  `CORE_XRM.usb_dn_en = $urandom;
	force  `CORE_XRM.usb_mode = $urandom;
	force  `CORE_XRM.usb_up_m_en = $urandom;
	force  `CORE_XRM.usb_up_p_en = $urandom;
	force  `CORE_XRM.utmi_suspend_n = $urandom;
	force  `CORE_XRM.utmifs_fs_edge_sel = $urandom;
	force  `CORE_XRM.utmifs_tx_dm = $urandom;
	force  `CORE_XRM.utmifs_tx_dp = $urandom;
	force  `CORE_XRM.utmifs_tx_enable_n = $urandom;
	force  `ANA_XRM.BB_ADC_I = $urandom;
	force  `ANA_XRM.BB_ADC_Q = $urandom;
	force  `ANA_XRM.BB_CLK_ADC_OUT = $urandom;
	force  `ANA_XRM.BB_RFINT = $urandom;
	force  `ANA_XRM.BB_RX_PKD_CLK = $urandom;
	force  `ANA_XRM.BB_RX_PKD_SAT = $urandom;
	force  `ANA_XRM.SPI_DO = $urandom;
	force  `ANA_XRM.utmifs_rx_dm = $urandom;
	force  `ANA_XRM.utmifs_rx_dp = $urandom;
	force  `ANA_XRM.utmifs_rx_rcv = $urandom;

 /*.scan_test_clock[[input]]*/          check_in_testmode (`ANA_XRM.scan_test_clock,`IOMUX_XRM.scan_test_clock,"");
 /*.test_en*/                           check_in_testmode (`QL_XRM.TEST_MODE_MBIST,`PAD_XRM.u_TEST_PAD.C,"TEST_MODE_MBIST");
 /*.sw_test_en*/                        check_in_testmode (`ANA_XRM.sw_test_en,`IOMUX_XRM.sw_test_en,"sw_test_en");
 /*.rf_test_en*/                        check_in_testmode (`ANA_XRM.rf_test_en,`IOMUX_XRM.rf_test_en,"rf_test_en");
 /*.bb_test_en*/                        check_in_testmode (`ANA_XRM.bb_test_en,`IOMUX_XRM.bb_test_en,"bb_test_en");
 /*.mbist_test_en*/                     check_in_testmode (`ANA_XRM.mbist_test_en,`IOMUX_XRM.mbist_test_en,"mbist_test_en");
 /*.bsd_test_en*/                       check_in_testmode (`ANA_XRM.bsd_test_en,`IOMUX_XRM.bsd_test_en,"bsd_test_en");
 /*.CLK_26M_OUT[[output]]*/             check_in_testmode (`IOMUX_XRM.osc_26m,`ANA_XRM.CLK_26M_OUT,"osc_26m");
 /*.CLK_26M[[input]]*/                  check_in_testmode (`QL_XRM.CLK_26M_RF,`CLK_XRM.clk_24m_rf,"CLK_26M_RF");
 /*.ADC_DATA[[output[10:0]]]*/          check_in_testmode (`SCUREG_XRM.ana_status1[31:21],`ANA_XRM.ADC_DATA[10:0],"ADC_DATA[10:0]");
 /*.ADC_VDET_INDEX[[output]]*/          check_in_testmode (`SCUREG_XRM.ana_status1[17],`ANA_XRM.ADC_VDET_INDEX,"ADC_VDET_INDEX");
 /*.DCDC_OCP_DET[[output]]*/            check_in_testmode (`IOMUX_XRM.dcdc_ocp_det,`ANA_XRM.DCDC_OCP_DET,"DCDC_OCP_DET");
 /*.DCDC_PWM_TEST[[output]]*/           check_in_testmode (`IOMUX_XRM.dcdc_pwm_test,`ANA_XRM.DCDC_PWM_TEST,"DCDC_PWM_TEST");
 /*.DCDC_START_TEST[[output]]*/         check_in_testmode (`IOMUX_XRM.dcdc_start_test,`ANA_XRM.DCDC_START_TEST,"DCDC_START_TEST");
 /*.DCDC_ZCD_TEST[[output]]*/           check_in_testmode (`IOMUX_XRM.dcdc_zcd_test,`ANA_XRM.DCDC_ZCD_TEST,"DCDC_ZCD_TEST");
 /*.DPLL_LOCK[[output]]*/               check_in_testmode (`IOMUX_XRM.dpll_lock,`ANA_XRM.DPLL_LOCK,"DPLL_LOCK");
 /*.DPLL_OUT_16M[[output]]*/            check_in_testmode (`CLK_XRM.pll_16m,`ANA_XRM.DPLL_OUT_16M,"DPLL_OUT_16M");
 /*.DPLL_OUT_24M[[output]]*/            check_in_testmode (`IOMUX_XRM.dpll_out_24m,`ANA_XRM.DPLL_OUT_24M,"DPLL_OUT_24M");
 /*.DPLL_OUT_192M[[output]]*/           check_in_testmode (`CLK_XRM.pll_192m,`ANA_XRM.DPLL_OUT_192M,"DPLL_OUT_192M");
 /*.DPLL_OUT_192M_TEST[[output]]*/      check_in_testmode (`IOMUX_XRM.dpll_out_192m_test,`ANA_XRM.DPLL_OUT_192M_TEST,"DPLL_OUT_192M_TEST");
 /*.LVD_BB[[output]]*/                  check_in_testmode (`SCU_XRM.lvd_bb,`ANA_XRM.LVD_BB,"LVD_BB");
 /*.POR_BB[[output]]*/                  check_in_testmode (`SCU_XRM.por_bb,`ANA_XRM.POR_BB,"POR_BB"); 
 /*.RCO32_CAL_CODE[[output[13:0]]]*/    check_in_testmode (`CORE_XRM.ana_status0[13:0],`ANA_XRM.RCO32_CAL_CODE[13:0],"RCO32_CAL_CODE[13:0]");                                               
 /*.RCO32_COARSE_DONE[[output]]*/       check_in_testmode (`IOMUX_XRM.rco32_coarse_done,`ANA_XRM.RCO32_COARSE_DONE,"RCO32_COARSE_DONE");      
 /*.RCO32_FINE_DONE[[output]]*/         check_in_testmode (`IOMUX_XRM.rco32_fine_done,`ANA_XRM.RCO32_FINE_DONE,"RCO32_FINE_DONE");                                               
 /*.RCO_32K_BB[[output]]*/              check_in_testmode (`CLK_XRM.rco_32k,`ANA_XRM.RCO_32K_BB,"RCO_32K_BB");                                               
 /*.ADC_CLK_SEL[[input[1:0]]]*/         check_in_testmode (`ANA_XRM.ADC_CLK_SEL[1:0],`SCU_XRM.ana_ctl4[11:10],"ADC_CLK_SEL[1:0]");                                               
 /*.ADC_GPIO33[[input[7:0]]]*/          check_in_testmode (`ANA_XRM.ADC_GPIO33[7:0],{4'b0,`PAD_XRM.ADC_IN[3:0]},"ADC_GPIO33[7:0]");                                               
 /*.ADC_GPIO_DIV[[input[1:0]]]*/        check_in_testmode (`ANA_XRM.ADC_GPIO_DIV[1:0],`SCU_XRM.ana_ctl3[5:4],"ADC_GPIO_DIV[1:0]");
 /*.ADC_GPIO_MUX[[input[2:0]]]*/        check_in_testmode (`ANA_XRM.ADC_GPIO_MUX[2:0],`SCU_XRM.ana_ctl3[8:6],"ADC_GPIO_MUX[2:0]");
 /*.ADC_INT_EN[[input]]*/               check_in_testmode (`ANA_XRM.ADC_INT_EN,`SCU_XRM.ana_ctl3[3],"ADC_INT_EN");
 /*.ADC_INT_MUX[[input[2:0]]]*/         check_in_testmode (`ANA_XRM.ADC_INT_MUX[2:0],`SCU_XRM.ana_ctl3[2:0],"ADC_INT_MUX[2:0]");
 /*.DCDC_LOGIC_MODE[[input]]*/          check_in_testmode (`ANA_XRM.DCDC_LOGIC_MODE,`SCU_XRM.ana_ctl4[2],"DCDC_LOGIC_MODE");
 /*.DCDC_RSV0[[input]]*/                check_in_testmode (`ANA_XRM.DCDC_RSV0,`SCU_XRM.ana_ctl4[1],"DCDC_RSV0");  
 /*.DCDC_RSV1[[input]]*/                check_in_testmode (`ANA_XRM.DCDC_RSV1,`SCU_XRM.ana_ctl4[0],"DCDC_RSV1");
 /*.ADC_START[[input]]*/                check_in_testmode (`ANA_XRM.ADC_START,`SCU_XRM.ana_ctl4[12],"ADC_START");
 /*.ADC_TEST_SEL[[input[1:0]]]*/        check_in_testmode (`ANA_XRM.ADC_TEST_SEL[1:0],`SCU_XRM.ana_ctl4[8:7],"ADC_TEST_SEL[1:0]");
 /*.ADC_VDET_BYPS[[input]]*/            check_in_testmode (`ANA_XRM.ADC_VDET_BYPS,`SCU_XRM.ana_ctl4[6],"ADC_VDET_BYPS");
 /*.BATDET_ADJ[[input[1:0]]]*/          check_in_testmode (`ANA_XRM.BATDET_ADJ[1:0],`SCU_XRM.ana_ctl4[14:13],"BATDET_ADJ[1:0]");
 /*.DCDC_FREQ_ADJ[[input[3:0]]]*/       check_in_testmode (`ANA_XRM.DCDC_FREQ_ADJ[3:0],`SCU_XRM.ana_ctl4[18:15],"DCDC_FREQ_ADJ[3:0]");
 /*.DCDC_OUT_ADJ[[input[1:0]]]*/        check_in_testmode (`ANA_XRM.DCDC_OUT_ADJ[1:0],`SCU_XRM.ana_ctl4[20:19],"DCDC_OUT_ADJ[1:0]");
 /*.DPLL_TEST_EN[[input]]*/             check_in_testmode (`ANA_XRM.DPLL_TEST_EN,`SCU_XRM.ana_ctl0[12],"DPLL_TEST_EN");
 /*.ENB_HV_LDO[[input]]*/               check_in_testmode (`ANA_XRM.ENB_HV_LDO,`SCU_XRM.ana_ctl0[31],"ENB_HV_LDO");
 /*.ENB_LDO_LP[[input]]*/               check_in_testmode (`ANA_XRM.ENB_LDO_LP,`SCU_XRM.ana_ctl0[29],"ENB_LDO_LP");
 /*.ENB_PMU_BG[[input]]*/               check_in_testmode (`ANA_XRM.ENB_PMU_BG,`SCU_XRM.ana_ctl0[30],"ENB_PMU_BG");
 /*.EN_ADC[[input]]*/                   check_in_testmode (`ANA_XRM.EN_ADC,`SCU_XRM.ana_ctl0[22],"EN_ADC");
 /*.EN_ADC_CNT_MODE[[input]]*/          check_in_testmode (`ANA_XRM.EN_ADC_CNT_MODE,`SCU_XRM.ana_ctl4[9],"EN_ADC_CNT_MODE");
 /*[[input[10:0]]].BB_DAC_I*/           check_in_testmode (`ANA_XRM.BB_DAC_I,`CORE_XRM.bb_dac_i[10:0],"BB_DAC_I");
 /*[[input[10:0]]].BB_DAC_Q*/           check_in_testmode (`ANA_XRM.BB_DAC_Q,`CORE_XRM.bb_dac_q[10:0],"BB_DAC_Q");
 /*[[input[10:0]]].BB_TX_GAIN*/         check_in_testmode (`ANA_XRM.BB_TX_GAIN,{~`CORE_XRM.bb_tx_gain[7:3], 3'h0, `CORE_XRM.bb_tx_gain[2:0]},"BB_TX_GAIN");
 /*[[input[13:0]]].RCO32_RCAL_EXT*/     check_in_testmode (`ANA_XRM.RCO32_RCAL_EXT,`SCUREG_XRM.ana_ctl2[29:16],"RCO32_RCAL_EXT");
 /*[[input[1:0]]].RCO32_CNT*/           check_in_testmode (`ANA_XRM.RCO32_CNT,`SCU_XRM.ana_ctl2[4:3],"RCO32_CNT");
 /*[[input[1:0]]].RCO32_TCAL*/          check_in_testmode (`ANA_XRM.RCO32_TCAL,`SCUREG_XRM.ana_ctl2[14:13],"RCO32_TCAL");
 /*[[input[1:0]]].VDT_BAT_ADJ*/         check_in_testmode (`ANA_XRM.VDT_BAT_ADJ,`SCU_XRM.ana_ctl3[28:27],"VDT_BAT_ADJ");
 /*[[input[2:0]]].HV_BG*/               check_in_testmode (`ANA_XRM.HV_BG,`SCU_XRM.ana_ctl1[18:16],"HV_BG");
 /*[[input[2:0]]].LDO_ADC_TRIM*/        check_in_testmode (`ANA_XRM.LDO_ADC_TRIM,`SCU_XRM.ana_ctl4[28:26],"LDO_ADC_TRIM");
 /*[[input[2:0]]].LDO_DG_TRIM*/         check_in_testmode (`ANA_XRM.LDO_DG_TRIM,`SCU_XRM.ana_ctl4[23:21],"LDO_DG_TRIM");
 /*[[input[2:0]]].LDO_LP_TRIM*/         check_in_testmode (`ANA_XRM.LDO_LP_TRIM,`SCU_XRM.ana_ctl3[31:29],"LDO_LP_TRIM");
 /*[[input[2:0]]].LDO_RF_TR*/           check_in_testmode (`ANA_XRM.LDO_RF_TR,`SCU_XRM.ana_ctl1[4:2],"LDO_RF_TR");
 /*[[input[2:0]]].LDO_XO_TRIM*/         check_in_testmode (`ANA_XRM.LDO_XO_TRIM,`SCU_XRM.ana_ctl4[31:29],"LDO_XO_TRIM");
 /*[[input[2:0]]].TEST_SEL*/            check_in_testmode (`ANA_XRM.TEST_SEL,`SCU_XRM.ana_ctl4[5:3],"TEST_SEL");
 /*[[input[3:0]]].LDO_LP_IBIAS_TRIM*/   check_in_testmode (`ANA_XRM.LDO_LP_IBIAS_TRIM,`SCU_XRM.ana_ctl3[26:23],"LDO_LP_IBIAS_TRIM");
 /*[[input[5:0]]].HV_LDO_TR*/           check_in_testmode (`ANA_XRM.HV_LDO_TR,`SCU_XRM.ana_ctl1[12:7],"HV_LDO_TR");
 /*[[input[6:0]]].BB_FREQ_HOP*/         check_in_testmode (`ANA_XRM.BB_FREQ_HOP,`CORE_XRM.bb_freq_hop[6:0],"BB_FREQ_HOP");
 /*[[input[7:0]]].BB_RX_AGC*/           check_in_testmode (`ANA_XRM.BB_RX_AGC,`CORE_XRM.bb_rx_agc[7:0],"BB_RX_AGC");
 /*[[input[7:0]]].BB_TEMP_COMP_TX_GAIN*/check_in_testmode (`ANA_XRM.BB_TEMP_COMP_TX_GAIN,`CORE_XRM.bb_temp_comp_tx_gain[7:0],"BB_TEMP_COMP_TX_GAIN");
 /*[[input]].BB_BT_RX_EN*/              check_in_testmode (`ANA_XRM.BB_BT_RX_EN,1'b0,"BB_BT_RX_EN");
 /*[[input]].BB_BT_SX_EN*/              check_in_testmode (`ANA_XRM.BB_BT_SX_EN,1'b0,"BB_BT_SX_EN");
 /*[[input]].BB_BT_TX_EN*/              check_in_testmode (`ANA_XRM.BB_BT_TX_EN,1'b0,"BB_BT_TX_EN");
 /*[[input]].BB_CLK_ADC_IN*/            check_in_testmode (`ANA_XRM.BB_CLK_ADC_IN,`CLK_XRM.rf_adc_clk,"BB_CLK_ADC_IN");
 /*[[input]].BB_CLK_DAC*/               check_in_testmode (`ANA_XRM.BB_CLK_DAC,`CLK_XRM.clk_48m_bb,"BB_CLK_DAC");
 /*[[input]].BB_DA_RX_PKD_RSTN*/        check_in_testmode (`ANA_XRM.BB_DA_RX_PKD_RSTN,`CORE_XRM.DA_RX_PKD_RSTN,"BB_DA_RX_PKD_RSTN");
 /*[[input]].CLK_26M_EN*/               check_in_testmode (`ANA_XRM.CLK_26M_EN,`SCU_XRM.ana_ctl0[4],"CLK_26M_EN");
 /*[[input]].CLK_EXT_IN*/               check_in_testmode (`ANA_XRM.CLK_EXT_IN,`IOMUX_XRM.clk_ext_in,"CLK_EXT_IN");
 /*[[input]].EN_32K_PAD*/               check_in_testmode (`ANA_XRM.EN_32K_PAD,`SCUREG_XRM.ana_ctl0[11],"EN_32K_PAD");
 /*[[input]].EN_BAT_DET*/               check_in_testmode (`ANA_XRM.EN_BAT_DET,`SCUREG_XRM.ana_ctl0[19],"EN_BAT_DET");
 /*[[input]].EN_CHIP_V33*/              check_in_testmode (`ANA_XRM.EN_CHIP_V33,`DUT_XRM.u_pad_ring.EN_CHIP_V33,"EN_CHIP_V33");
 /*[[input]].EN_DCDC*/                  check_in_testmode (`ANA_XRM.EN_DCDC,`SCUREG_XRM.ana_ctl0[28],"EN_DCDC");
 /*[[input]].EN_DCDC_OCP*/              check_in_testmode (`ANA_XRM.EN_DCDC_OCP,`SCUREG_XRM.ana_ctl0[15],"EN_DCDC_OCP");
 /*[[input]].EN_DCDC_TEST*/             check_in_testmode (`ANA_XRM.EN_DCDC_TEST,`SCUREG_XRM.ana_ctl0[14],"EN_DCDC_TEST");
 /*[[input]].EN_DCDC_VDT*/              check_in_testmode (`ANA_XRM.EN_DCDC_VDT,`SCUREG_XRM.ana_ctl0[17],"EN_DCDC_VDT");
 /*[[input]].EN_DPLL*/                  check_in_testmode (`ANA_XRM.EN_DPLL,`CLK_XRM.mux_dpll_sel,"EN_DPLL");
 /*[[input]].EN_DPLL_LOCK_BYPS*/        check_in_testmode (`ANA_XRM.EN_DPLL_LOCK_BYPS,`SCUREG_XRM.ana_ctl0[13],"EN_DPLL_LOCK_BYPS");
 /*[[input]].EN_LDO_ADC*/               check_in_testmode (`ANA_XRM.EN_LDO_ADC,`SCUREG_XRM.ana_ctl0[25],"EN_LDO_ADC");
 /*[[input]].EN_LDO_RF*/                check_in_testmode (`ANA_XRM.EN_LDO_RF,`SCUREG_XRM.ana_ctl0[27],"EN_LDO_RF");
 /*[[input]].EN_LDO_XO*/                check_in_testmode (`ANA_XRM.EN_LDO_XO,`CLK_XRM.mux_ldoxo_sel,"EN_LDO_XO");
 /*[[input]].EN_RCO32K_BIAS*/           check_in_testmode (`ANA_XRM.EN_RCO32K_BIAS,`SCUREG_XRM.ana_ctl1[23],"EN_RCO32K_BIAS");
 /*[[input]].EN_RCO_32K*/               check_in_testmode (`ANA_XRM.EN_RCO_32K,`SCUREG_XRM.ana_ctl0[21],"EN_RCO_32K");
 /*[[input]].EN_VDT_BAT*/               check_in_testmode (`ANA_XRM.EN_VDT_BAT,`SCUREG_XRM.ana_ctl0[18],"EN_VDT_BAT");
 /*[[input]].EN_VDT_RF*/                check_in_testmode (`ANA_XRM.EN_VDT_RF,`SCUREG_XRM.ana_ctl0[16],"EN_VDT_RF");
 /*[[input]].HV_BAT_BYPASS*/            check_in_testmode (`ANA_XRM.HV_BAT_BYPASS,`SCUREG_XRM.ana_ctl1[5],"HV_BAT_BYPASS");
 /*[[input]].HV_LDO_LOAD*/              check_in_testmode (`ANA_XRM.HV_LDO_LOAD,`SCUREG_XRM.ana_ctl1[6],"HV_LDO_LOAD");
 /*[[input]].HV_LDO_USB_BAT*/           check_in_testmode (`ANA_XRM.HV_LDO_USB_BAT,`SCUREG_XRM.ana_ctl1[15],"HV_LDO_USB_BAT");
 /*[[input]].LDO_RF_BYPASS*/            check_in_testmode (`ANA_XRM.LDO_RF_BYPASS,`SCUREG_XRM.ana_ctl1[0],"LDO_RF_BYPASS");
 /*[[input]].LDO_RF_LOAD*/              check_in_testmode (`ANA_XRM.LDO_RF_LOAD,`SCUREG_XRM.ana_ctl1[1],"LDO_RF_LOAD");
 /*[[input]].RCO32_BIAS_ADJ*/           check_in_testmode (`ANA_XRM.RCO32_BIAS_ADJ,`SCUREG_XRM.ana_ctl1[22],"RCO32_BIAS_ADJ");
 /*[[input]].RCO32_COARSE_CAL_EN*/      check_in_testmode (`ANA_XRM.RCO32_COARSE_CAL_EN,`SCUREG_XRM.ana_ctl2[31],"RCO32_COARSE_CAL_EN");
 /*[[input]].RCO32_FINE_CAL_EN*/        check_in_testmode (`ANA_XRM.RCO32_FINE_CAL_EN,`SCUREG_XRM.ana_ctl2[30],"RCO32_FINE_CAL_EN");
 /*[[input]].RCO32_FOUT*/               check_in_testmode (`ANA_XRM.RCO32_FOUT,`SCUREG_XRM.ana_ctl2[15],"RCO32_FOUT");
 /*[[input]].RCO32_RCAL_EXTEN*/         check_in_testmode (`ANA_XRM.RCO32_RCAL_EXTEN,`SCUREG_XRM.ana_ctl2[12],"RCO32_RCAL_EXTEN");
 /*[[input]].RESETN_RF*/                check_in_testmode (`ANA_XRM.RESETN_RF,`IOMUX_XRM.resetn_rf,"RESETN_RF");
 /*[[input]].SPI_CLK*/                  check_in_testmode (`ANA_XRM.SPI_CLK,`IOMUX_XRM.rf_spis_clk_ana,"SPI_CLK");
 /*[[input]].SPI_CSN*/                  check_in_testmode (`ANA_XRM.SPI_CSN,`IOMUX_XRM.rf_spis_csn_ana,"SPI_CSN");
 /*[[input]].SPI_DI*/                   check_in_testmode (`ANA_XRM.SPI_DI,`IOMUX_XRM.rf_spis_mosi_ana,"SPI_DI");
 /*[[input]].usb_dn_en*/                check_in_testmode (`ANA_XRM.usb_dn_en,`CORE_XRM.usb_dn_en,"usb_dn_en");
 /*[[input]].usb_mode*/                 check_in_testmode (`ANA_XRM.usb_mode,`CORE_XRM.usb_mode,"usb_mode");
 /*[[input]].usb_up_m_en*/              check_in_testmode (`ANA_XRM.usb_up_m_en,`CORE_XRM.usb_up_m_en,"usb_up_m_en");
 /*[[input]].usb_up_p_en*/              check_in_testmode (`ANA_XRM.usb_up_p_en,`CORE_XRM.usb_up_p_en,"usb_up_p_en");
 /*[[input]].utmi_suspend_n*/           check_in_testmode (`ANA_XRM.utmi_suspend_n,`CORE_XRM.utmi_suspend_n,"utmi_suspend_n");
 /*[[input]].utmifs_fs_edge_sel*/       check_in_testmode (`ANA_XRM.utmifs_fs_edge_sel,`CORE_XRM.utmifs_fs_edge_sel,"utmifs_fs_edge_sel");
 /*[[input]].utmifs_tx_dm*/             check_in_testmode (`ANA_XRM.utmifs_tx_dm,`CORE_XRM.utmifs_tx_dm,"utmifs_tx_dm");
 /*[[input]].utmifs_tx_dp*/             check_in_testmode (`ANA_XRM.utmifs_tx_dp,`CORE_XRM.utmifs_tx_dp,"utmifs_tx_dp");
 /*[[input]].utmifs_tx_enable_n*/       check_in_testmode (`ANA_XRM.utmifs_tx_enable_n,`CORE_XRM.utmifs_tx_enable_n,"utmifs_tx_enable_n");
 /*[[output[9:0]]].BB_ADC_I*/           check_in_testmode (`BB_XRM.rxdata_i[9:0],`ANA_XRM.BB_ADC_I,"BB_ADC_I");
 /*[[output[9:0]]].BB_ADC_Q*/           check_in_testmode (`BB_XRM.rxdata_q[9:0],`ANA_XRM.BB_ADC_Q,"BB_ADC_Q");
 /*[[output]].BB_CLK_ADC_OUT*/          check_in_testmode (`BB_XRM.clk_bt_adc,`ANA_XRM.BB_CLK_ADC_OUT,"BB_CLK_ADC_OUT");
 /*[[output]].BB_RFINT*/                check_in_testmode (`CORE_XRM.rf_int,`ANA_XRM.BB_RFINT,"BB_RFINT");
 /*[[output]].BB_RX_PKD_CLK*/           check_in_testmode (`DUT_XRM.bb_rx_pkd_clk,`ANA_XRM.BB_RX_PKD_CLK,"BB_RX_PKD_CLK");
 /*[[output]].BB_RX_PKD_SAT*/           check_in_testmode (`CORE_XRM.bb_rx_pkd_sat,`ANA_XRM.BB_RX_PKD_SAT,"BB_RX_PKD_SAT");
 /*[[output]].SPI_DO*/                  check_in_testmode (`IOMUX_XRM.rf_spis_miso_ana,`ANA_XRM.SPI_DO,"SPI_DO");
 /*[[output]].utmifs_rx_dm*/            check_in_testmode (`USBPHY_XRM.U_DWC_otg_piu.utmifs_rx_dm,`ANA_XRM.utmifs_rx_dm,"utmifs_rx_dm");
 /*[[output]].utmifs_rx_dp*/            check_in_testmode (`USBPHY_XRM.U_DWC_otg_piu.utmifs_rx_dp,`ANA_XRM.utmifs_rx_dp,"utmifs_rx_dp");
 /*[[output]].utmifs_rx_rcv*/           check_in_testmode (`USBPHY_XRM.U_DWC_otg_piu.utmifs_rx_rcv,`ANA_XRM.utmifs_rx_rcv,"utmifs_rx_rcv");
        $display("CLK_SDC_CYCLE The %d times loop", i);
  end // for

  if (!error_count == 0) 
	$display ("CNT test FAIL, error_count = %d",error_count);
    else
        $display("CNT test succeessfully ");
endtask: ana_connect_dig


// check task 
task check_in_testmode (left_sigin,right_sigal,string name); 
//  #10;// it would tested the value of singal 10ns ago;
  if (left_sigin !== right_sigal) 
    begin
      error_count = error_count + 1;
      $display("%t %s left signal is %b, right signal is %b test FAIL!!!!!!!!!!",$realtime,name,left_sigin,right_sigal);
    end //else
    //$display("%t %s left signal is %b, right signal is %b test RIGHT",$realtime,name,left_sigin,right_sigal);
  #10;
endtask: check_in_testmode

