`timescale 1ns/1ps

module user_def;
	defparam  u_spi_flash0.Init_File = "./inputs/soc_top/sim/tests/s_1_002_scu_remap_flash/flash.hex";
endmodule
