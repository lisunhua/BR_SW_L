`timescale 1ns/1ps


module user_def;
	defparam CLT.m_uart.Input_Udata = "./inputs/soc_top/sim/tests/d_1_24E_bb_rom_cmd_sleep_hw_roc_32k_wp_gpio/uart_clt.cm";
	defparam SVR.m_uart.Input_Udata = "./inputs/soc_top/sim/tests/d_1_24E_bb_rom_cmd_sleep_hw_roc_32k_wp_gpio/uart_svr.cm";
endmodule
