`timescale 1ns/1ps


module user_def;
	defparam CLT.m_uart.Input_Udata = "./inputs/soc_top/sim/tests/d_1_252_bb_rom_cmd_sleep_sw_roc_32k/uart_clt.cm";
	defparam SVR.m_uart.Input_Udata = "./inputs/soc_top/sim/tests/d_1_252_bb_rom_cmd_sleep_sw_roc_32k/uart_svr.cm";
endmodule
