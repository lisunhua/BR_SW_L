`timescale 1ns/1ps

module user_def;
	defparam  soc_tb.u_spi_flash0.Init_File = "./inputs/soc_top/sim/tests/s_1_007_scu_scan_xip_flash/flash.hex";
endmodule
