`timescale 1ns/1ps


module user_def;
	defparam CLT.m_uart.Input_Udata = "./inputs/soc_top/sim/tests/d_1_24F_bb_rom_cmd_sleep_hw_osc_32k/uart_clt.cm";
	defparam SVR.m_uart.Input_Udata = "./inputs/soc_top/sim/tests/d_1_24F_bb_rom_cmd_sleep_hw_osc_32k/uart_svr.cm";
endmodule
