`timescale 1ns/1ps

module user_def;
	defparam soc_tb.m_uart.Input_Udata = "./inputs/soc_top/sim/tests/s_1_657_scu_change_pclk_async_uart0_rx/uart.cm";
endmodule
