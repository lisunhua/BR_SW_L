`timescale 1ns/1ps


module user_def;
	defparam CLT.m_uart.Input_Udata = "./inputs/soc_top/sim/tests/d_1_24D_bb_rom_cmd_sleep_hw_osc_24m_div_32k_baud_1800/uart_clt.cm";
	defparam SVR.m_uart.Input_Udata = "./inputs/soc_top/sim/tests/d_1_24D_bb_rom_cmd_sleep_hw_osc_24m_div_32k_baud_1800/uart_svr.cm";
endmodule
