`timescale 1ns/1ps

module user_def;
	defparam soc_tb.u_usb_host_sim.DATA_PATH = "./inputs/soc_top/sim/tests/s_1_251_bb_rom_usb_sacn/usb_host_sim_data.txt";
endmodule
